aser